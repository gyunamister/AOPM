DEFINE  "c1: An order must be delivered in 200"  AS
ENTITY "Order"
ASSOCIATE "Order", "Item", "Package", "Route"
VALIDATE "membership", IN, {"Gold"}
EVALUATE "Throughput", <, 200;

DEFINE  "c2: An availability of item must be checked before picking"  AS
ENTITY "Item"
VALIDATE "pick_item", IN, {activity}
EVALUATE "check_availability", EVENTUALLY, "pick_item";