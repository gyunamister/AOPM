DEFINE "cf1"  AS
CONTEXT "omap"={"Order":{"foreach"}}
FILTER "event"
EVALUATE "Throughput", <, 72; 